magic
tech scmos
timestamp 1554908150
use __CIF2__  __CIF2___0
timestamp 1554908150
transform 1 0 0 0 1 0
box 0 0 5000 5000
<< end >>
